class transaction;
  rand bit [7:0]data;
  rand bit rd_wr;
  bit mosi;
  bit miso;
  
endclass
